module Segment_Display_7(
    input [3:0] valor , // Número 0 -> 9
    output reg [6:0]hex // (a,b,c,d,e,g,h)
);

    always @(*) begin
        case (valor)

           4'd0: hex = 7'b1000000; // 0
           4'd1: hex = 7'b1111001; // 1
           4'd2: hex = 7'b0100100; // 2
           4'd3: hex = 7'b0110000; // 3
           4'd4: hex = 7'b0011001; // 4
           4'd5: hex = 7'b0010010; // 5
           4'd6: hex = 7'b0000010; // 6
           4'd7: hex = 7'b1111000; // 7
           4'd8: hex = 7'b0000000; // 8
           4'd9: hex = 7'b0010000; // 9

           default: hex = 7'b1111111;
        endcase
    end
endmodule
