module Freq_Div_1Hz (
    input clk,          
    output reg tick_1s  
);

    reg [25:0] contador;
    
    // Frequência FPGA: 50MHz
    always @(posedge clk) begin
        if (contador == 50000000 - 1) begin
            contador <= 0;
            tick_1s <= 1; // Ativa o pulso
            
        end else begin
            contador <= contador + 1;
            tick_1s <= 0; // Desativa o pulso
        end
    end
endmodule
